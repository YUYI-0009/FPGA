module mux3_1(
input wire [1:0] s,
input wire [7:0] a,b,c,
output reg [7:0] y
);
always @(s) begin
	if(s==2'b10) y=c;
	else if(s==2'b01) y=b;
	else y=a;
	end
endmodule