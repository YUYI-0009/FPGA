module mux3_1(
	input wire [7:0] a,b,c,
	input wire [1:0] s,
	output reg [7:0] y
);
always @(s,a,b,c) begin
	if(s==2'b00) y=a;
	else if(s==2'b01) y=b;
	else if(s==2'b10) y=c;
	else y=a;
	end
endmodule 
