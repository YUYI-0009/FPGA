module mux2_1(
	input wire [7:0] a,b,
	input wire s,
	output reg [7:0] y
);
 always @(s,a,b) begin
	if(s==1'b0) y=a;
	else y=b;
	end
endmodule
	